00
FF
00
E0
22
30
6E
00
6D
01
FD
15
A2
50
FE
1E
F1
65
A2
4A
D0
11
C0
7F
C1
3F
D0
11
A2
50
FE
1E
F1
55
7E
02
4E
3C
6E
00
F0
07
30
00
12
28
12
0A
6E
00
62
02
C0
7F
C1
3F
A2
50
FE
1E
F1
55
A2
4A
D0
11
7E
02
3E
3C
12
34
00
EE
80
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
00
