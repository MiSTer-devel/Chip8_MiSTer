00
FF
00
E0
00
FE
60
00
61
00
62
00
63
00
64
00
65
00
66
00
67
00
68
00
69
00
6A
00
6B
00
6C
00
6D
00
6E
00
6F
00
F0
15
F0
18
A0
00
12
00
